module MUL(
        clk,
        rst_n,
        a,
        B,
        result
        );

    input [31:0] A,B;
    output reg [63:0] result;

    wire [31:0] pp [0:31]; 
    wire [63:0] sum, carry;
    wire [63:0] final_sum;
    //===================================================//
    d32_d28 L1 (
        .clk(clk),
        .rst_n(rst_n),
        .pp(pp), 
        .s1(s1),
        .c1(c1),
        .pp1(pp1)
    );

    d28_d19 L2 (
        .clk(clk),
        .rst_n(rst_n),
        .pp1(pp1), 
        .s1(s1),
        .c1(c1),
        .s2(s2),
        .c2(c2),
        .pp2(pp2),
        .remain2(remain2)
    );

    d19_d13 L3 (
        .clk(clk),
        .rst_n(rst_n),
        .pp2(pp2), 
        .remain2(remain2),
        .s2(s2),
        .c2(c2),
        .s3(s3),
        .c3(c3),
        .pp3(pp3),
        .remain3(remain3)
    );

    //===================================================//


    genvar i;
    generate
        for (i = 0; i < 32; i = i+1) begin : gen_pp
            assign pp[i] = A & {32{B[i]}};
        end
    endgenerate
    
    assign result = sum + carry;


endmodule 


module HA (
    input  a,
    input  b,
    output sum,
    output carry
    );

    assign sum   = a ^ b;
    assign carry = a & b;
endmodule

module FA (
    input  a,
    input  b,
    input  cin,
    output sum,
    output cout
    );

    assign sum  = a ^ b ^ cin;
    assign cout = (a & b) | (b & cin) | (a & cin);

endmodule

module d32_d28 (
    clk,
    rst_n,
    pp,
    s1,
    c1,
    pp1
    );

    input clk, rst_n;
    input [31:0] pp [0:31];
    output reg [19:0] s1;
    output reg [19:0] c1;
    output reg [31:0] pp1 [0:31];

    wire [19:0] s;
    wire [19:0] c;
    //--------------------------//
    // [28]
    HA ha0 (pp[28][0], pp[27][1], s[0], c[0]);
    //[29]
    FA fa0 (pp[29][0], pp[28][1], pp[27][2], s[1], c[1]);
    HA ha1 (pp[26][3], pp[25][4], s[2], c[2]);
    // [30]
    FA fa1 (pp[30][0], pp[29][1], pp[28][2], s[3], c[3]);
    FA fa2 (pp[27][3], pp[26][4], pp[25][5], s[4], c[4]);
    HA ha2 (pp[24][6], pp[23][7], s[5], c[5]);
    // [31]
    FA fa3 (pp[31][0], pp[30][1], pp[29][2], s[6], c[6]);
    FA fa4 (pp[28][3], pp[27][4], pp[26][5], s[7], c[7]);
    FA fa5 (pp[25][6], pp[24][7], pp[23][8], s[8], c[8]);
    HA ha3 (pp[22][9], pp[21][10], s[9], c[9]);
    // [30]
    FA fa6 (pp[30][2], pp[29][3], pp[28][4], s[10], c[10]);
    FA fa7 (pp[27][5], pp[26][6], pp[25][7], s[11], c[11]);
    FA fa8 (pp[24][8], pp[23][9], pp[22][10], s[12], c[12]);
    HA ha4 (pp[21][11], pp[20][12], s[13], c[13]);
    // [29]
    FA fa9  (pp[29][4], pp[28][5], pp[27][6], s[14], c[14]);
    FA fa10 (pp[26][7], pp[25][8], pp[24][9], s[15], c[15]);
    FA fa11 (pp[23][10], pp[22][11], pp[21][12], s[16], c[16]);
    //[28]
    FA fa12 (pp[28][6], pp[27][7], pp[26][8], s[17], c[17]);
    FA fa13 (pp[25][9], pp[24][10], pp[23][11], s[18], c[18]);
    //[27]
    FA fa14 (pp[27][8], pp[26][9], pp[25][10], s[19], c[19]);

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            s1 <= 20'd0;
            c1 <= 20'd0;
        end 
        else begin
            s1 <= s;
            c1 <= c;
            pp1 <= pp;
        end
    end


endmodule

module d28_d19 (
    clk,
    rst_n,
    pp1
    s1,
    c1,
    s2,
    c2,
    pp2,
    remain2
    );

    input clk, rst_n;
    input [31:0] pp1 [0:31];
    input [19:0] s1;
    input [19:0] c1;
    output reg [161:0] s2, C2;
    output reg [31:0] pp2 [0:31];
    output reg [8:0] remain2;

    wire [161:0] s, c;
//---------------------------------------//
    //19
    HA ha1 (pp1[19][0], pp1[18][1], s[0], c[0]);
    //20
    FA fa1 (pp1[20][0], pp1[19][1], pp1[18][2], s[1], c[1]);
    HA ha2 (pp1[17][3], pp1[16][4], s[2], c[2]);
    //21
    FA fa2 (pp1[21][0], pp1[20][1], pp1[19][2], s[3], c[3]);
    FA fa3 (pp1[18][3], pp1[17][4], pp1[16][5], s[4], c[4]);
    HA ha3 (pp1[15][6], pp1[14][7], s[5], c[5]);
    //22
    FA fa4 (pp1[22][0], pp1[21][1], pp1[20][2], s[6], c[6]);
    FA fa5 (pp1[19][3], pp1[18][4], pp1[17][5], s[7], c[7]);
    FA fa6 (pp1[16][6], pp1[15][7], pp1[14][8], s[8], c[8]);
    HA ha4 (pp1[13][9], pp1[12][10], s[9], c[9]);
    //23
    FA fa7 (pp1[23][0], pp1[22][1], pp1[21][2], s[10], c[10]);
    FA fa8 (pp1[20][3], pp1[19][4], pp1[18][5], s[11], c[11]);
    FA fa9 (pp1[17][6], pp1[16][7], pp1[15][8], s[12], c[12]);
    FA fa10 (pp1[14][9], pp1[13][10], pp1[12][11], s[13], c[13]);
    HA ha5 (pp1[11][12], pp1[10][13], s[14], c[14]);   
    //24
    FA fa11 (pp1[24][0], pp1[23][1], pp1[22][2], s[15], c[15]);
    FA fa12 (pp1[21][3], pp1[20][4], pp1[19][5], s[16], c[16]);
    FA fa13 (pp1[18][6], pp1[17][7], pp1[16][8], s[17], c[17]);
    FA fa14 (pp1[15][9], pp1[14][10], pp1[13][11], s[18], c[18]);
    FA fa15 (pp1[12][12], pp1[11][13], pp1[10][14], s[19], c[19]);    
    HA ha6 (pp1[9][15], pp1[8][16], s[20], c[20]);    
    //25
    FA fa16 (pp1[25][0], pp1[24][1], pp1[23][2], s[21], c[21]);
    FA fa17 (pp1[22][3], pp1[21][4], pp1[20][5], s[22], c[22]);
    FA fa18 (pp1[19][6], pp1[18][7], pp1[17][8], s[23], c[23]);
    FA fa19 (pp1[16][9], pp1[15][10], pp1[14][11], s[24], c[24]);
    FA fa20 (pp1[13][12], pp1[12][13], pp1[11][14], s[25], c[25]); 
    FA fa21 (pp1[10][15], pp1[9][16], pp1[8][17], s[26], c[26]);    
    HA ha7 (pp1[7][18], pp1[6][19], s[27], c[27]); 
    //26
    FA fa22 (pp1[26][0], pp1[25][1], pp1[24][2], s[28], c[28]);
    FA fa23 (pp1[23][3], pp1[22][4], pp1[21][5], s[29], c[29]);
    FA fa24 (pp1[20][6], pp1[19][7], pp1[18][8], s[30], c[30]);
    FA fa25 (pp1[17][9], pp1[16][10], pp1[15][11], s[31], c[31]);
    FA fa26 (pp1[14][12], pp1[13][13], pp1[12][14], s[32], c[32]); 
    FA fa27 (pp1[11][15], pp1[10][16], pp1[9][17], s[33], c[33]);    
    FA fa28 (pp1[8][18], pp1[7][19], pp1[6][20], s[34], c[34]); 
    HA ha8 (pp1[5][21], pp1[4][22], s[35], c[35]); 
    //27
    FA fa29 (pp1[27][0], pp1[26][1], pp1[25][2], s[36], c[36]);
    FA fa30 (pp1[24][3], pp1[23][4], pp1[22][5], s[37], c[37]);
    FA fa31 (pp1[21][6], pp1[20][7], pp1[19][8], s[38], c[38]);
    FA fa32 (pp1[18][9], pp1[17][10], pp1[16][11], s[39], c[39]);
    FA fa33 (pp1[15][12], pp1[14][13], pp1[13][14], s[40], c[40]); 
    FA fa34 (pp1[12][15], pp1[11][16], pp1[10][17], s[41], c[41]);    
    FA fa35 (pp1[9][18], pp1[8][19], pp1[7][20], s[42], c[42]); 
    FA fa37 (pp1[6][21], pp1[5][22], pp1[4][23], s[43], c[43]); 
    HA ha9 (pp1[3][24], pp1[2][25], s[44], c[44]);  
    //28[27][1]
    FA fa38 (pp1[26][2], pp1[25][3], pp1[24][4], s[45], c[45]);
    FA fa39 (pp1[23][5], pp1[22][6], pp1[21][7], s[46], c[46]);
    FA fa40 (pp1[20][8], pp1[19][9], pp1[18][10], s[47], c[47]);
    FA fa41 (pp1[17][11], pp1[16][12], pp1[15][13], s[48], c[48]);
    FA fa42 (pp1[14][14], pp1[13][15], pp1[12][16], s[49], c[49]); 
    FA fa43 (pp1[11][17], pp1[10][18], pp1[19][19], s[50], c[50]);    
    FA fa44 (pp1[8][20], pp1[7][21], pp1[6][22], s[51], c[51]); 
    FA fa45 (pp1[5][23], pp1[4][24], pp1[3][25], s[52], c[52]); 
    FA fa46 (pp1[2][26], pp1[1][27], pp1[0][28], s[53], c[53]);  
    //29[25][4]
    FA fa47 (pp1[24][5], pp1[23][6], pp1[22][7], s[54], c[54]);
    FA fa48 (pp1[21][8], pp1[20][9], pp1[19][10], s[55], c[55]);
    FA fa49 (pp1[18][11], pp1[17][12], pp1[16][13], s[56], c[56]);
    FA fa50 (pp1[15][14], pp1[14][15], pp1[13][16], s[57], c[57]);
    FA fa51 (pp1[12][17], pp1[11][18], pp1[10][19], s[58], c[58]); 
    FA fa52 (pp1[9][20], pp1[8][21], pp1[7][22], s[59], c[59]);    
    FA fa53 (pp1[6][23], pp1[5][24], pp1[4][25], s[60], c[60]); 
    FA fa54 (pp1[3][26], pp1[2][27], pp1[1][28], s[61], c[61]); 
    FA fa55 (pp1[0][29], s1[1], s1[2], s[62], c[62]); 
    //30[23][7]
    FA fa56 (pp1[22][8], pp1[21][9], pp1[20][10], s[63], c[63]);
    FA fa57 (pp1[19][11], pp1[18][12], pp1[17][13], s[64], c[64]);
    FA fa58 (pp1[16][14], pp1[15][15], pp1[14][16], s[65], c[65]);
    FA fa59 (pp1[13][17], pp1[12][18], pp1[11][19], s[66], c[66]);
    FA fa60 (pp1[10][20], pp1[9][21], pp1[8][22], s[67], c[67]); 
    FA fa61 (pp1[7][23], pp1[6][24], pp1[5][25], s[68], c[68]);    
    FA fa62 (pp1[4][26], pp1[3][27], pp1[2][28], s[69], c[69]); 
    FA fa63 (pp1[1][29], pp1[0][30], s1[3], s[70], c[70]); 
    FA fa64 (s1[4], s1[5], c1[1], s[71], c[71]); 
    //31[21][10]
    FA fa65 (pp1[20][11], pp1[19][12], pp1[18][13], s[72], c[72]);
    FA fa66 (pp1[17][14], pp1[16][15], pp1[15][16], s[73], c[73]);
    FA fa67 (pp1[14][17], pp1[13][18], pp1[12][19], s[74], c[74]);
    FA fa68 (pp1[11][20], pp1[10][21], pp1[9][22], s[75], c[75]);
    FA fa69 (pp1[8][23], pp1[7][24], pp1[6][25], s[76], c[76]); 
    FA fa70 (pp1[5][26], pp1[4][27], pp1[3][28], s[77], c[77]);    
    FA fa71 (pp1[2][29], pp1[1][30], pp1[0][31], s[78], c[78]); 
    FA fa72 (s1[6], s1[7], s1[8], s[79], c[79]); 
    FA fa73 (s1[9], c1[3], c1[4], s[80], c[80]); 
    //30[20][12]+1
    FA fa74 (pp1[19][13], pp1[18][14], pp1[17][15], s[81], c[81]);
    FA fa75 (pp1[16][16], pp1[15][17], pp1[14][18], s[82], c[82]);
    FA fa76 (pp1[13][19], pp1[12][20], pp1[11][21], s[83], c[83]);
    FA fa77 (pp1[10][22], pp1[9][23], pp1[8][24], s[84], c[84]);
    FA fa78 (pp1[7][25], pp1[6][26], pp1[5][27], s[85], c[85]); 
    FA fa79 (pp1[4][28], pp1[3][29], pp1[2][30], s[86], c[86]);    
    FA fa80 (pp1[1][31], pp1[31][1], s1[10], s[87], c[87]); 
    FA fa81 (s1[11], s1[12], s1[13], s[88], c[88]); 
    FA fa82 (c1[6], c1[7], c1[8], s[89], c[89]); 
    //29[21][12]+2
    FA fa83 (pp1[20][13], pp1[19][14], pp1[18][15], s[90], c[90]);
    FA fa84 (pp1[17][16], pp1[16][17], pp1[15][18], s[91], c[91]);
    FA fa85 (pp1[14][19], pp1[13][20], pp1[12][21], s[92], c[92]);
    FA fa86 (pp1[11][22], pp1[10][23], pp1[9][24], s[93], c[93]);
    FA fa87 (pp1[8][25], pp1[7][26], pp1[6][27], s[94], c[94]); 
    FA fa88 (pp1[5][28], pp1[4][29], pp1[3][30], s[95], c[95]);    
    FA fa89 (pp1[2][31], pp1[31][2], pp1[30][3], s[96], c[96]); 
    FA fa90 (s1[14], s1[15], s1[16], s[97], c[97]); 
    FA fa91 (c1[10], c1[11], c1[12], s[98], c[98]); 
    //28[23][11]+3
    FA fa92 (pp1[22][12], pp1[21][13], pp1[20][14], s[99], c[99]);
    FA fa93 (pp1[19][15], pp1[18][16], pp1[17][17], s[100], c[100]);
    FA fa94 (pp1[16][18], pp1[15][19], pp1[14][20], s[101], c[101]);
    FA fa95 (pp1[13][21], pp1[12][22], pp1[11][23], s[102], c[102]);
    FA fa96 (pp1[10][24], pp1[9][25], pp1[8][26], s[103], c[103]); 
    FA fa97 (pp1[7][27], pp1[6][28], pp1[5][29], s[104], c[104]);    
    FA fa98 (pp1[4][30], pp1[3][31], pp1[31][3], s[105], c[105]); 
    FA fa99 (pp1[30][4], pp1[29][5], s1[17], s[106], c[106]); 
    FA fa100 (s1[18], c1[14], c1[15], s[107], c[107]); 
    //27[25][10]+4
    FA fa101 (pp1[24][11], pp1[23][12], pp1[22][13], s[108], c[108]);
    FA fa102 (pp1[21][14], pp1[20][15], pp1[19][16], s[109], c[109]);
    FA fa103 (pp1[18][17], pp1[17][18], pp1[16][19], s[110], c[110]);
    FA fa104 (pp1[15][20], pp1[14][21], pp1[13][22], s[111], c[111]);
    FA fa105 (pp1[12][23], pp1[11][24], pp1[10][25], s[112], c[112]); 
    FA fa106 (pp1[9][26], pp1[8][27], pp1[7][28], s[113], c[113]);    
    FA fa107 (pp1[6][29], pp1[5][30], pp1[4][31], s[114], c[114]); 
    FA fa108 (pp1[31][4], pp1[30][5], pp1[29][6], s[115], c[115]); 
    FA fa109 (pp1[28][7], s1[19], c1[17], s[116], c[116]); 
    // 26+5
    FA fa110 (pp1[26][10], pp1[25][11], pp1[24][12], s[117], c[117]);
    FA fa111 (pp1[23][13], pp1[22][14], pp1[21][15], s[118], c[118]);
    FA fa112 (pp1[20][16], pp1[19][17], pp1[18][18], s[119], c[119]);
    FA fa113 (pp1[17][19], pp1[16][20], pp1[15][21], s[120], c[120]);
    FA fa114 (pp1[14][22], pp1[13][23], pp1[12][24], s[121], c[121]); 
    FA fa115 (pp1[11][25], pp1[10][26], pp1[9][27], s[122], c[122]);    
    FA fa116 (pp1[8][28], pp1[7][29], pp1[6][30], s[123], c[123]); 
    FA fa117 (pp1[5][31], pp1[31][5], pp1[30][6], s[124], c[124]); 
    FA fa118 (pp1[29][7], pp1[28][8], pp1[27][9], s[125], c[125]); 
    //25+6
    FA fa119 (pp1[25][12], pp1[24][13], pp1[23][14], s[126], c[126]);
    FA fa120 (pp1[22][15], pp1[21][16], pp1[20][17], s[127], c[127]);
    FA fa121 (pp1[19][18], pp1[18][19], pp1[17][20], s[128], c[128]);
    FA fa122 (pp1[16][21], pp1[15][22], pp1[14][23], s[129], c[129]);
    FA fa123 (pp1[13][24], pp1[12][25], pp1[11][26], s[130], c[130]);
    FA fa124 (pp1[10][27], pp1[9][28], pp1[8][29], s[131], c[131]);
    FA fa125 (pp1[7][30], pp1[6][31], pp1[31][6], s[132], c[132]);
    FA fa126 (pp1[30][7], pp1[29][8], pp1[28][9], s[133], c[133]);
    // 24+7
    FA fa127 (pp1[24][14], pp1[23][15], pp1[22][16], s[134], c[134]);
    FA fa128 (pp1[21][17], pp1[20][18], pp1[19][19], s[135], c[135]);
    FA fa129 (pp1[18][20], pp1[17][21], pp1[16][22], s[136], c[136]);
    FA fa130 (pp1[15][23], pp1[14][24], pp1[13][25], s[137], c[137]);
    FA fa131 (pp1[12][26], pp1[11][27], pp1[10][28], s[138], c[138]);
    FA fa132 (pp1[9][29], pp1[8][30], pp1[7][31], s[139], c[139]);
    FA fa133 (pp1[31][7], pp1[30][8], pp1[29][9], s[140], c[140]);
    // 23+8
    FA fa134 (pp1[23][16], pp1[22][17], pp1[21][18], s[141], c[141]);
    FA fa135 (pp1[20][19], pp1[19][20], pp1[18][21], s[142], c[142]);
    FA fa136 (pp1[17][22], pp1[16][23], pp1[15][24], s[143], c[143]);
    FA fa137 (pp1[14][25], pp1[13][26], pp1[12][27], s[144], c[144]);
    FA fa138 (pp1[11][28], pp1[10][29], pp1[9][30], s[145], c[145]);
    FA fa139 (pp1[8][31], pp1[31][8], pp1[30][9], s[146], c[146]);
    // 22+9
    FA fa140 (pp1[22][18], pp1[21][19], pp1[20][20], s[147], c[147]);
    FA fa141 (pp1[19][21], pp1[18][22], pp1[17][23], s[148], c[148]);
    FA fa142 (pp1[16][24], pp1[15][25], pp1[14][26], s[149], c[149]);
    FA fa143 (pp1[13][27], pp1[12][28], pp1[11][29], s[150], c[150]);
    FA fa144 (pp1[10][30], pp1[9][31], pp1[31][9], s[151], c[151]);
    // 21+10
    FA fa145 (pp1[21][20], pp1[20][21], pp1[19][22], s[152], c[152]);
    FA fa146 (pp1[18][23], pp1[17][24], pp1[16][25], s[153], c[153]);
    FA fa147 (pp1[15][26], pp1[14][27], pp1[13][28], s[154], c[154]);
    FA fa148 (pp1[12][29], pp1[11][30], pp1[10][31], s[155], c[155]);
    // 20+11
    FA fa149 (pp1[20][22], pp1[19][23], pp1[18][24], s[156], c[156]);
    FA fa150 (pp1[17][25], pp1[16][26], pp1[15][27], s[157], c[157]);
    FA fa151 (pp1[14][28], pp1[13][29], pp1[12][30], s[158], c[158]);
    // 19+12
    FA fa152 (pp1[19][24], pp1[18][25], pp1[17][26], s[159], c[159]);
    FA fa153 (pp1[16][27], pp1[15][28], pp1[14][29], s[160], c[160]);
    // 18+13
    FA fa154 (pp1[18][26], pp1[17][27], pp1[16][28], s[161], c[161]);

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            s2 <= 162'd0;
            c2 <= 162'd0;
            remain2 <= 9'd0;
        end 
        else begin
            s2 <= s;
            c2 <= c;
            pp2 <= pp1;
            remain2 <= {c1[19], c1[17], c1[16], c1[13], c1[9], c1[5], c1[2], c1[0], s1[0]};
        end
    end

endmodule

module d19_d13 (
    clk,
    rst_n,
    pp2
    remain2,
    s2,
    c2,
    s3,
    c3,
    pp3,
    remain3
    );

    input clk, rst_n;
    input [31:0] pp2 [0:31];
    input [155:0] s2, C2;
    input [8:0] remain2;
    output reg [197:0] s3, c3;
    output reg [31:0] pp3 [0:31];
    output reg [17:0] remain3;

    wire [197:0] s, c;
//------------------------------//
    // 13
    HA ha1 (pp2[13][0], pp2[12][1], s[0], c[0]);
    // 14
    FA fa1 (pp2[14][0], pp2[13][1], pp2[12][2], s[1], c[1]);
    HA ha2 (pp2[11][3], pp2[10][4], s[2], c[2]);
    // 15
    FA fa2 (pp2[15][0], pp2[14][1], pp2[13][2], s[3], c[3]);
    FA fa3 (pp2[12][3], pp2[11][4], pp2[10][5], s[4], c[4]);
    HA ha3 (pp2[9][6], pp2[8][7], s[5], c[5]);
    // 16
    FA fa4 (pp2[16][0], pp2[15][1], pp2[14][2], s[6], c[6]);
    FA fa5 (pp2[13][3], pp2[12][4], pp2[11][5], s[7], c[7]);
    FA fa6 (pp2[10][6], pp2[9][7], pp2[8][8], s[8], c[8]);
    HA ha4 (pp2[7][9], pp2[6][10], s[9], c[9]);
    // 17
    FA fa7 (pp2[17][0], pp2[16][1], pp2[15][2], s[10], c[10]);
    FA fa8 (pp2[14][3], pp2[13][4], pp2[12][5], s[11], c[11]);
    FA fa9 (pp2[11][6], pp2[10][7], pp2[9][8], s[12], c[12]);
    FA fa10 (pp2[8][9], pp2[7][10], pp2[6][11], s[13], c[13]);
    HA ha5 (pp2[5][12], pp2[4][13], s[14], c[14]); 
    // 18
    FA fa11 (pp2[18][0], pp2[17][1], pp2[16][2], s[15], c[15]);
    FA fa12 (pp2[15][3], pp2[14][4], pp2[13][5], s[16], c[16]);
    FA fa13 (pp2[12][6], pp2[11][7], pp2[10][8], s[17], c[17]);
    FA fa14 (pp2[9][9], pp2[8][10], pp2[7][11], s[18], c[18]);
    FA fa15 (pp2[6][12], pp2[5][13], pp2[4][14], s[19], c[19]);    
    HA ha6 (pp2[3][15], pp2[2][16], s[20], c[20]); 
    // 19[18][1]
    FA fa16 (pp2[17][2], pp2[16][3], pp2[15][4], s[21], c[21]);
    FA fa17 (pp2[14][5], pp2[13][6], pp2[12][7], s[22], c[22]);
    FA fa18 (pp2[11][8], pp2[10][9], pp2[9][10], s[23], c[23]);
    FA fa19 (pp2[8][11], pp2[7][12], pp2[6][13], s[24], c[24]);
    FA fa20 (pp2[5][14], pp2[4][15], pp2[3][16], s[25], c[25]); 
    FA fa21 (pp2[2][17], pp2[1][18], pp2[0][19], s[26], c[26]); 
    // 20[16][4]
    FA fa22 (pp2[15][5], pp2[14][6], pp2[13][7], s[27], c[27]);
    FA fa23 (pp2[12][8], pp2[11][9], pp2[10][10], s[28], c[28]);
    FA fa24 (pp2[9][11], pp2[8][12], pp2[7][13], s[29], c[29]);
    FA fa25 (pp2[6][14], pp2[5][15], pp2[4][16], s[30], c[30]);
    FA fa26 (pp2[3][17], pp2[2][18], pp2[1][19], s[31], c[31]); 
    FA fa27 (pp2[0][20], s2[1], s2[2], s[32], c[32]);     
    // 21[14][7]
    FA fa28 (pp2[13][8], pp2[12][9], pp2[11][10], s[33], c[33]);
    FA fa29 (pp2[10][11], pp2[9][12], pp2[8][13], s[34], c[34]);
    FA fa30 (pp2[7][14], pp2[6][15], pp2[5][16], s[35], c[35]);
    FA fa31 (pp2[4][17], pp2[3][18], pp2[2][19], s[36], c[36]);
    FA fa32 (pp2[1][20], pp2[0][21], s2[3], s[37], c[37]); 
    FA fa33 (s2[4], s2[5], c2[1], s[38], c[38]);
    // 22[12][10]
    FA fa34 (pp2[11][11], pp2[10][12], pp2[9][13], s[39], c[39]);
    FA fa35 (pp2[8][14], pp2[7][15], pp2[6][16], s[40], c[40]);
    FA fa36 (pp2[5][17], pp2[4][18], pp2[3][19], s[41], c[41]);
    FA fa37 (pp2[2][20], pp2[1][21], pp2[0][22], s[42], c[42]);
    FA fa38 (s2[6], s2[7], s2[8], s[43], c[43]);
    FA fa39 (s2[9], c2[3], c2[4], s[44], c[44]);
    // 23[10][13]
    FA fa40 (pp2[9][14], pp2[8][15], pp2[7][16], s[45], c[45]);
    FA fa41 (pp2[6][17], pp2[5][18], pp2[4][19], s[46], c[46]);
    FA fa42 (pp2[3][20], pp2[2][21], pp2[1][22], s[47], c[47]);
    FA fa43 (pp2[0][23], s2[10], s2[11], s[48], c[48]);
    FA fa44 (s2[12], s2[13], s2[14], s[49], c[49]);
    FA fa45 (c2[6], c2[7], c2[8], s[50], c[50]);
    // 24[8][16]
    FA fa46 (pp2[7][17], pp2[6][18], pp2[5][19], s[51], c[51]);
    FA fa47 (pp2[4][20], pp2[3][21], pp2[2][22], s[52], c[52]);
    FA fa48 (pp2[1][23], pp2[0][24], s2[15], s[53], c[53]);
    FA fa49 (s2[16], s2[17], s2[18], s[54], c[54]);
    FA fa50 (s2[19], s2[20], c2[10], s[55], c[55]);
    FA fa51 (c2[11], c2[12], c2[13], s[56], c[56]);
    // 25[6][19]
    FA fa52 (pp2[5][20], pp2[4][21], pp2[3][22], s[57], c[57]);
    FA fa53 (pp2[2][23], pp2[1][24], pp2[0][25], s[58], c[58]);
    FA fa54 (s2[21], s2[22], s2[23], s[59], c[59]);
    FA fa55 (s2[24], s2[25], s2[26], s[60], c[60]);
    FA fa56 (s2[27], c2[15], c2[16], s[61], c[61]);
    FA fa57 (c2[17], c2[18], c2[19], s[62], c[62]);
    // 26[4][22]
    FA fa58 (pp2[3][23], pp2[2][24], pp2[1][25], s[63], c[63]);
    FA fa59 (pp2[0][26], s2[28], s2[29], s[64], c[64]);
    FA fa60 (s2[30], s2[31], s2[32], s[65], c[65]);
    FA fa61 (s2[33], s2[34], s2[35], s[66], c[66]);
    FA fa62 (c2[21], c2[22], c2[23], s[67], c[67]);
    FA fa63 (c2[24], c2[25], c2[26], s[68], c[68]);
    // 27[2][25]
    FA fa64 (pp2[1][26], pp2[0][27], s2[36], s[69], c[69]);
    FA fa65 (s2[37], s2[38], s2[39], s[70], c[70]);
    FA fa66 (s2[40], s2[41], s2[42], s[71], c[71]);
    FA fa67 (s2[43], s2[44], c2[28], s[72], c[72]);
    FA fa68 (c2[29], c2[30], c2[31], s[73], c[73]);
    FA fa69 (c2[32], c2[33], c2[34], s[74], c[74]);
    // 28
    FA fa70 (remain2[0], s2[45], s2[46], s[75], c[75]);
    FA fa71 (s2[47], s2[48], s2[49], s[76], c[76]);
    FA fa72 (s2[50], s2[51], s2[52], s[77], c[77]);
    FA fa73 (s2[53], c2[36], c2[37], s[78], c[78]);
    FA fa74 (c2[38], c2[39], c2[40], s[79], c[79]);
    FA fa75 (c2[41], c2[42], c2[43], s[80], c[80]);
    // 29
    FA fa76 (remain2[1], s2[54], s2[55], s[81], c[81]);
    FA fa77 (s2[56], s2[57], s2[58], s[82], c[82]);
    FA fa78 (s2[59], s2[60], s2[61], s[83], c[83]);
    FA fa79 (s2[62], c2[45], c2[46], s[84], c[84]);
    FA fa80 (c2[47], c2[48], c2[49], s[85], c[85]);
    FA fa81 (c2[50], c2[51], c2[52], s[86], c[86]);
    // 30
    FA fa82 (remain2[2], s2[63], s2[64], s[87], c[87]);
    FA fa83 (s2[65], s2[66], s2[67], s[88], c[88]);
    FA fa84 (s2[68], s2[69], s2[70], s[89], c[89]);
    FA fa85 (s2[71], c2[54], c2[55], s[90], c[90]);
    FA fa86 (c2[56], c2[57], c2[58], s[91], c[91]);
    FA fa87 (c2[59], c2[60], c2[61], s[92], c[92]);
    // 31
    FA fa88 (remain2[3], s2[72], s2[73], s[93], c[93]);
    FA fa89 (s2[74], s2[75], s2[76], s[94], c[94]);
    FA fa90 (s2[77], s2[78], s2[79], s[95], c[95]);
    FA fa91 (s2[80], c2[63], c2[64], s[96], c[96]);
    FA fa92 (c2[65], c2[66], c2[67], s[97], c[97]);
    FA fa93 (c2[68], c2[69], c2[70], s[98], c[98]);
    // 30
    FA fa94 (remain2[4], s2[81], s2[82], s[99], c[99]);
    FA fa95 (s2[83], s2[84], s2[85], s[100], c[100]);
    FA fa96 (s2[86], s2[87], s2[88], s[101], c[101]);
    FA fa97 (s2[89], c2[72], c2[73], s[102], c[102]);  
    FA fa98 (c2[74], c2[75], c2[76], s[103], c[103]);
    FA fa99 (c2[77], c2[78], c2[79], s[104], c[104]);
    // 29
    FA fa100 (remain2[5], s2[90], s2[91], s[105], c[105]);
    FA fa101 (s2[92], s2[93], s2[94], s[106], c[106]);
    FA fa102 (s2[95], s2[96], s2[97], s[107], c[107]);
    FA fa103 (s2[98], c2[81], c2[82], s[108], c[108]);
    FA fa104 (c2[83], c2[84], c2[85], s[109], c[109]);
    FA fa105 (c2[86], c2[87], c2[88], s[110], c[110]);
    // 28
    FA fa106 (remain2[6], s2[99], s2[100], s[111], c[111]);
    FA fa107 (s2[101], s2[102], s2[103], s[112], c[112]);
    FA fa108 (s2[104], s2[105], s2[106], s[113], c[113]);
    FA fa109 (s2[107], c2[90], c2[91], s[114], c[114]);
    FA fa110 (c2[92], c2[93], c2[94], s[115], c[115]);
    FA fa111 (c2[95], c2[96], c2[97], s[116], c[116]);
    // 27
    FA fa112 (remain2[7], s2[108], s2[109], s[117], c[117]);
    FA fa113 (s2[110], s2[111], s2[112], s[118], c[118]);
    FA fa114 (s2[113], s2[114], s2[115], s[119], c[119]);
    FA fa115 (s2[116], c2[99], c2[100], s[120], c[120]);
    FA fa116 (c2[101], c2[102], c2[103], s[121], c[121]);
    FA fa117 (c2[104], c2[105], c2[106], s[122], c[122]);
    // 26
    FA fa118 (remain2[8], s2[117], s2[118], s[123], c[123]);
    FA fa119 (s2[119], s2[120], s2[121], s[124], c[124]);
    FA fa120 (s2[122], s2[123], s2[124], s[125], c[125]);
    FA fa121 (s2[125], c2[108], c2[109], s[126], c[126]);
    FA fa122 (c2[110], c2[111], c2[112], s[127], c[127]);
    FA fa123 (c2[113], c2[114], c2[115], s[128], c[128]);
    // 25[28][9]+6
    FA fa124 (pp2[27][10], s2[126], s2[127], s[129], c[129]);
    FA fa125 (s2[128], s2[129], s2[130], s[130], c[130]);
    FA fa126 (s2[131], s2[132], s2[133], s[131], c[131]);
    FA fa127 (c2[117], c2[118], c2[119], s[132], c[132]);
    FA fa128 (c2[120], c2[121], c2[122], s[133], c[133]);
    FA fa129 (c2[123], c2[124], c2[125], s[134], c[134]);
    // 24[29][9]+7
    FA fa130 (s2[134], s2[135], s2[136], s[135], c[135]);
    FA fa131 (s2[137], s2[138], s2[139], s[136], c[136]);
    FA fa132 (s2[140], c2[126], c2[127], s[137], c[137]);
    FA fa133 (c2[128], c2[129], c2[130], s[138], c[138]);
    FA fa134 (c2[131], c2[132], c2[133], s[139], c[139]);
    FA fa135 (pp2[28][10], pp2[27][11], pp2[26][12], s[140], c[140]);
    // 23[30][9]+8
    FA fa136 (s2[141], s2[142], s2[143], s[141], c[141]);
    FA fa137 (s2[144], s2[145], s2[146], s[142], c[142]);
    FA fa138 (c2[134], c2[135], c2[136], s[143], c[143]);
    FA fa139 (c2[137], c2[138], c2[139], s[144], c[144]);
    FA fa140 (c2[140], pp2[29][10], pp2[28][11], s[145], c[145]);
    FA fa141 (pp2[27][12], pp2[26][13], pp2[25][14], s[146], c[146]);
    // 22[31][9]+9
    FA fa142 (s2[147], s2[148], s2[149], s[147], c[147]);
    FA fa143 (s2[150], s2[151], c2[141], s[148], c[148]);
    FA fa144 (c2[142], c2[143], c2[144], s[149], c[149]);
    FA fa145 (c2[145], c2[146], pp2[30][10], s[150], c[150]);
    FA fa146 (pp2[29][11], pp2[28][12], pp2[27][13], s[151], c[151]);
    FA fa147 (pp2[26][14], pp2[25][15], pp2[24][16], s[152], c[152]);
    // 21[10][31]+10
    FA fa148 (s2[152], s2[153], s2[154], s[153], c[153]);
    FA fa149 (s2[155], c2[147], c2[148], s[154], c[154]);
    FA fa150 (c2[149], c2[150], c2[151], s[155], c[155]);
    FA fa151 (pp2[31][10], pp2[30][11], pp2[29][12], s[156], c[156]);
    FA fa152 (pp2[28][13], pp2[27][14], pp2[26][15], s[157], c[157]);
    FA fa153 (pp2[25][16], pp2[24][17], pp2[23][18], s[158], c[158]);
    // 20[12][30]+11
    FA fa154 (s2[156], s2[157], s2[158], s[159], c[159]);
    FA fa155 (c2[152], c2[153], c2[154], s[160], c[160]);
    FA fa156 (c2[155], pp2[11][31], pp2[31][11], s[161], c[161]);
    FA fa157 (pp2[30][12], pp2[29][13], pp2[28][14], s[162], c[162]);
    FA fa158 (pp2[27][15], pp2[26][16], pp2[25][17], s[163], c[163]);
    FA fa159 (pp2[24][18], pp2[23][19], pp2[22][20], s[164], c[164]);
    // 19[14][29]+12
    FA fa160 (s2[159], s2[160], c2[156], s[165], c[165]);
    FA fa161 (c2[157], c2[158], pp2[13][30], s[166], c[166]);
    FA fa162 (pp2[12][31], pp2[31][12], pp2[30][13], s[167], c[167]);
    FA fa163 (pp2[29][14], pp2[28][15], pp2[27][16], s[168], c[168]);
    FA fa164 (pp2[26][17], pp2[25][18], pp2[24][19], s[169], c[169]);
    FA fa165 (pp2[23][20], pp2[22][21], pp2[21][22], s[170], c[170]);
    //18[16][28]+13
    FA fa166 (s2[161], c2[159], c2[160], s[171], c[171]);
    FA fa167 (pp2[15][29], pp2[14][30], pp2[13][31], s[172], c[172]);
    FA fa168 (pp2[31][13], pp2[30][14], pp2[29][15], s[173], c[173]);
    FA fa169 (pp2[28][16], pp2[27][17], pp2[26][18], s[174], c[174]);
    FA fa170 (pp2[25][19], pp2[24][20], pp2[23][21], s[175], c[175]);
    FA fa171 (pp2[22][22], pp2[21][23], pp2[20][24], s[176], c[176]);
    // 17+14
    FA fa172 (pp2[17][28], pp2[16][29], pp2[15][30], s[177], c[177]);
    FA fa173 (pp2[14][31], pp2[31][14], c2[161], s[178], c[178]);
    FA fa174 (pp2[30][15], pp2[29][16], pp2[28][17], s[179], c[179]);
    FA fa175 (pp2[27][18], pp2[26][19], pp2[25][20], s[180], c[180]);
    FA fa176 (pp2[24][21], pp2[23][22], pp2[22][23], s[181], c[181]);
    FA fa177 (pp2[21][24], pp2[20][25], pp2[19][26], s[182], c[182]);
    // 16+15
    FA fa178 (pp2[16][30], pp2[15][31], pp2[31][15], s[183], c[183]);
    FA fa179 (pp2[30][16], pp2[29][17], pp2[28][18], s[184], c[184]);
    FA fa180 (pp2[27][19], pp2[26][20], pp2[25][21], s[185], c[185]);
    FA fa181 (pp2[24][22], pp2[23][23], pp2[22][24], s[186], c[186]);
    FA fa182 (pp2[21][25], pp2[20][26], pp2[19][27], s[187], c[187]);
    // 15+16
    FA fa183 (pp2[16][31], pp2[31][16], pp2[30][17], s[188], c[188]);
    FA fa184 (pp2[29][18], pp2[28][19], pp2[27][20], s[189], c[189]);
    FA fa185 (pp2[26][21], pp2[25][22], pp2[24][23], s[190], c[190]);
    FA fa186 (pp2[23][24], pp2[22][25], pp2[21][26], s[191], c[191]);
    // 14+15
    FA fa187 (pp2[31][17], pp2[30][18], pp2[29][19], s[192], c[192]);
    FA fa188 (pp2[28][20], pp2[27][21], pp2[26][22], s[193], c[193]);
    FA fa189 (pp2[25][23], pp2[24][24], pp2[23][25], s[194], c[194]);
    // 13+14
    FA fa190 (pp2[31][18], pp2[30][19], pp2[29][20], s[195], c[195]);
    FA fa191 (pp2[28][21], pp2[27][22], pp2[26][23], s[196], c[196]);
    // 12+15
    FA fa192 (pp2[31][19], pp2[30][20], pp2[29][21], s[197], c[197]);

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            s3 <= 198'd0;
            c3 <= 198'd0;
            remain2 <= 9'd0;
        end 
        else begin
            s3 <= s;
            c3 <= c;
            pp3 <= pp2;
            remain3 <= {c2[116], c2[107], c2[98], c2[89], c2[80], 
                    c2[71], c2[62], c2[53], c2[44], c2[35], c2[27], 
                    c2[20], c2[14], c2[9], c2[5], c2[2], c2[0], remain2[0]};
        end
    end

endmodule